* My First Circuit

V1 1 0 DC 5V
R1 1 2 1k
R2 2 0 1k

.DC V1 0 5 0.1
.PRINT DC V(2)

.END
